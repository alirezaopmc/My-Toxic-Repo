library verilog;
use verilog.vl_types.all;
entity ArrayMultiplier_6x6_TB is
    generic(
        N               : integer := 6;
        M               : integer := 6
    );
end ArrayMultiplier_6x6_TB;
