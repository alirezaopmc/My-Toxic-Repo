library verilog;
use verilog.vl_types.all;
entity SixteenBitAdderTest is
end SixteenBitAdderTest;
