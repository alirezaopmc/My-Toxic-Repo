library verilog;
use verilog.vl_types.all;
entity bcd_test is
end bcd_test;
