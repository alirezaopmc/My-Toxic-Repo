library verilog;
use verilog.vl_types.all;
entity TestHalfAdder is
end TestHalfAdder;
