library verilog;
use verilog.vl_types.all;
entity TestFullAdder is
end TestFullAdder;
