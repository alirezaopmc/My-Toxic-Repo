library verilog;
use verilog.vl_types.all;
entity CarrySelectAdder_16bit_3_3_6_4_TB is
    generic(
        N               : integer := 16
    );
end CarrySelectAdder_16bit_3_3_6_4_TB;
