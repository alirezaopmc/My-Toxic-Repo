library verilog;
use verilog.vl_types.all;
entity FourBitAdderTest is
end FourBitAdderTest;
